----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 02/18/2021 08:31:47 PM
-- Design Name: 
-- Module Name: debounce - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity debounce is
    Port ( clk : in STD_LOGIC;
           btn : in STD_LOGIC;
           dbnc : out STD_LOGIC);
end debounce;

architecture Behavioral of debounce is
signal sreg : std_logic_vector(1 downto 0);
signal samples: std_logic_vector(2 downto 0); --max samples: 4
signal counter: std_logic_vector(26 downto 0);

begin
    process(clk)
        begin
            if (rising_edge(clk)) then
                if (unsigned(counter) < 124999999) then
                    counter <= std_logic_vector(unsigned(counter) + 1);
                else
                    counter <= (others => '0');            
                end if;
                sreg(1) <= sreg(0);
                sreg(0) <= btn;
                if (sreg(1) = '1') then
                    if(unsigned(samples) < 4) then
                        samples <= std_logic_vector(unsigned(samples) + 1);
                    end if;
                else
                    samples <= (others => '0');
                end if;
                if (unsigned(samples) = 4) then
                    dbnc <= '1';
                else
                    dbnc <= '0';
                end if;            
           end if;
   end process;

end Behavioral;
